module consts

pub const sampling_rate = 44100
